----------------------------------------------------------------------------------
-- Company:        ITESM - CQ
-- Engineer:       Rick
-- 
-- Create Date:    10:19:48 11/08/2017 
-- Design Name: 
-- Module Name:    VGA_DISPLAY - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description:    Here a drawing will be created 
--  
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
-- Commonly used libraries
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

entity VGA_DISPLAY is
  Generic
	 ( n : integer := 14;   -- Number of Address bus lines, for an image of 128x128 pixels
	   m : integer := 8);   -- Number of Data bus lines
  port (
	 Xin       : in  STD_LOGIC_VECTOR(9 downto 0); -- Column screen coordinate
	 Yin       : in  STD_LOGIC_VECTOR(9 downto 0); -- Row screen coordinate
	 En        : in  STD_LOGIC; -- When '1', pixels can be drawn 
	 Enable60  : in STD_LOGIC; --Enable for duck
	 Enable2   : in STD_LOGIC; --Enable for strawberry
	 Enable3   : in STD_LOGIC; --Enable for anviel
	 rightB    : in STD_LOGIC; --Right button
	 leftB     : in STD_LOGIC; --Left button
	 rst       : in STD_LOGIC; --Reset
	 clk       : in STD_LOGIC; --Clock from FPGA
	 FlagOut   : out STD_LOGIC; --Tells the score when to count
	 R   		  : out STD_LOGIC_VECTOR(2 downto 0); -- 3-bit Red channel
	 G   		  : out STD_LOGIC_VECTOR(2 downto 0); -- 3-bit Green channel
	 B   		  : out STD_LOGIC_VECTOR(1 downto 0));-- 2-bit Blue channel
end VGA_DISPLAY;


architecture Behavioral of VGA_DISPLAY is
  -- Embedded signal to group the colors into 1-byte
  -- The colors will be as follows:
  --  R2 R1 R0 G2 G1 G0 B1 B0
  signal Color : STD_LOGIC_VECTOR(7 downto 0); 
  --Addresses for the different images that will be displayed
  signal AddressChar : STD_LOGIC_VECTOR(n-1 downto 0); --Duck
  signal AddressObj  : STD_LOGIC_VECTOR(n-3 downto 0); --Strawberry
  signal AddressObj2 : STD_LOGIC_VECTOR(n-3 downto 0); --Anviel
  signal AddressKok : STD_LOGIC_VECTOR(n-7 downto 0); --Heart
  signal AddressGO : STD_LOGIC_VECTOR(n-1 downto 0); --Pantalla Game Over
  signal AddressBS : STD_LOGIC_VECTOR(n-1 downto 0); --Pantalla de Inicio

  signal Data:    STD_LOGIC_VECTOR(m-1 downto 0);
  
  --Types of roms that will be used
  type objectImage is array (0 to (64**2) - 1) of STD_LOGIC_VECTOR (7 downto 0);
  type characterImage is array (0 to (128**2) - 1) of STD_LOGIC_VECTOR (7 downto 0);
  type kokoroImage is array (0 to (2**8) - 1) of STD_LOGIC_VECTOR (7 downto 0); --n=8 (8 bits) porque 2^n=2^8=256
  type GO_Screen is array (0 to (2**14) - 1) of STD_LOGIC_VECTOR (7 downto 0);
  type Begin_Screen is array (0 to (2**14) - 1) of STD_LOGIC_VECTOR (7 downto 0);
 
 
  constant ImageBS : Begin_Screen := (
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"4C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",
x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",
x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",
x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",
x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",
x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",
x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",
x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",
x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",
x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",
x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",
x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",
x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",
x"8C",x"8C",x"8C",x"8C",x"8C",x"8C",x"4C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F9",x"F9",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FF",x"FF",x"F5",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FA",x"FF",x"F5",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F9",x"F5",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FF",x"FF",x"F9",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"90",x"FA",x"FA",x"F9",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FA",x"FF",x"FA",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F5",x"FF",x"FF",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FA",x"FF",x"F9",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"51",x"FF",x"FF",x"FF",x"FF",x"FA",x"F4",x"F4",
x"F4",x"F4",x"F9",x"FF",x"FA",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"FA",x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"FF",x"FF",x"F5",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FA",x"FF",x"FA",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"4D",
x"FF",x"FF",x"F5",x"F4",x"FF",x"FF",x"F4",x"F4",
x"F4",x"F4",x"F5",x"FF",x"FA",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F5",x"FF",x"FF",x"F9",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FA",x"FF",x"F9",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"DB",
x"FF",x"B5",x"F4",x"F4",x"FA",x"FF",x"F4",x"F4",
x"F4",x"F4",x"F5",x"FF",x"FE",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"FF",x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FA",x"FF",x"F5",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"71",x"FF",
x"B6",x"8C",x"F4",x"F4",x"FA",x"FE",x"F4",x"F4",
x"F4",x"F4",x"F4",x"FF",x"FE",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FA",x"FF",x"FF",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F9",x"FA",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F9",x"FA",x"F5",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F5",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F5",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F5",x"D6",x"BA",
x"96",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"DB",x"FF",
x"2C",x"8C",x"F4",x"F4",x"F5",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FF",x"FF",x"FF",x"FA",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F5",
x"FF",x"FF",x"FF",x"FF",x"F4",x"F4",x"F4",x"FA",
x"FF",x"FF",x"FF",x"FA",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FF",x"FF",x"FF",x"FF",
x"F5",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",x"F9",x"FA",
x"F4",x"F4",x"F9",x"F4",x"F4",x"F4",x"F4",x"FF",
x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"FA",x"F9",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F5",x"FF",x"FF",x"FF",x"FF",
x"FF",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"4D",x"FF",x"BA",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",
x"F5",x"FF",x"FA",x"F4",x"FF",x"FF",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F9",x"FF",
x"FF",x"F4",x"F9",x"FF",x"F9",x"F4",x"F4",x"F5",
x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F5",x"FF",x"FF",x"F5",x"F5",x"FF",
x"FA",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"FF",x"FF",x"F5",x"F9",x"FA",x"FF",x"FF",x"FF",
x"F5",x"F5",x"FF",x"FA",x"F4",x"F4",x"F4",x"FF",
x"FF",x"F5",x"F4",x"F4",x"F4",x"FF",x"FF",x"FF",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FA",x"FF",x"FF",x"F5",x"90",x"2C",
x"2C",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"96",x"FF",x"71",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",
x"FF",x"FF",x"F4",x"F4",x"FA",x"FF",x"F5",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F9",x"FF",x"FE",
x"F4",x"F4",x"F5",x"FF",x"F5",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FF",x"F5",x"F5",x"FA",x"FF",x"FF",
x"FE",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F5",x"FF",x"FF",x"F4",x"F4",x"F4",x"FF",
x"FA",x"F4",x"F4",x"F4",x"F4",x"F5",x"FA",x"FE",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"FA",x"F5",
x"F4",x"F5",x"FF",x"FF",x"F4",x"F4",x"F4",x"FA",
x"FF",x"F9",x"F4",x"F4",x"FA",x"FF",x"F9",x"FF",
x"F9",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FF",x"FA",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"DB",x"FF",x"2C",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"FA",
x"FF",x"F5",x"F4",x"F4",x"F9",x"FF",x"F9",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F5",x"FF",x"FF",x"F4",
x"F4",x"F4",x"F9",x"FF",x"FE",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FF",x"F5",x"F4",x"F4",x"F4",x"F5",
x"FF",x"FF",x"FA",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",x"FF",
x"FF",x"F4",x"F5",x"FF",x"FF",x"FF",x"FF",x"FE",
x"FF",x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",x"FA",
x"FF",x"F9",x"F4",x"F4",x"FF",x"F9",x"F4",x"FF",
x"FA",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"2C",x"FF",x"DF",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"FF",
x"FF",x"F4",x"F4",x"F4",x"F5",x"FF",x"F9",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",
x"F4",x"F4",x"FF",x"FF",x"FF",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FF",x"FA",x"F4",x"F4",x"F4",x"F4",
x"FF",x"FF",x"F5",x"F4",x"F4",x"F4",x"FA",x"FF",
x"FF",x"F4",x"F4",x"F5",x"F5",x"F4",x"F4",x"F4",
x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",x"F9",
x"FF",x"FA",x"F4",x"FA",x"FF",x"F4",x"F4",x"FF",
x"FA",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"FF",x"FF",x"F9",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"4D",x"FF",x"BA",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"FF",x"FF",x"F4",x"FA",x"FF",
x"F5",x"F4",x"F4",x"F4",x"F5",x"FF",x"FA",x"F4",
x"F4",x"F4",x"F4",x"FF",x"FF",x"F5",x"F4",x"F4",
x"F4",x"FA",x"FF",x"FF",x"FF",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",x"FA",
x"FF",x"FA",x"F4",x"F4",x"F4",x"F5",x"FF",x"FF",
x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FF",x"FE",x"F4",x"F4",x"F4",x"F9",
x"FF",x"FA",x"F4",x"FF",x"FA",x"F4",x"F4",x"FF",
x"FE",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FE",x"FF",x"FF",x"FF",x"DA",x"71",
x"2C",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"71",x"FF",x"96",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"FF",x"FF",x"F4",x"FF",x"FF",
x"F4",x"F4",x"F4",x"F4",x"F5",x"FF",x"FA",x"F4",
x"F4",x"F4",x"F9",x"FF",x"FA",x"F4",x"F4",x"F4",
x"F5",x"FF",x"FA",x"FF",x"FF",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",x"FF",
x"FF",x"F4",x"F4",x"F4",x"F4",x"FF",x"FF",x"FA",
x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",x"F5",
x"FF",x"FA",x"F9",x"FF",x"F4",x"F4",x"F4",x"FF",
x"FE",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F9",x"FA",x"FF",x"FF",
x"FF",x"BA",x"4D",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"71",x"FF",x"96",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"FF",x"F4",x"FF",x"FF",x"F9",x"FF",x"F9",
x"F4",x"F4",x"F4",x"F4",x"F5",x"FF",x"FA",x"F4",
x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",
x"FF",x"FF",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",
x"F5",x"FF",x"FF",x"FA",x"F4",x"F4",x"FE",x"FF",
x"F5",x"F4",x"F4",x"F4",x"FA",x"FF",x"F4",x"FA",
x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"FE",x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",
x"FF",x"FE",x"FF",x"FA",x"F4",x"F4",x"F4",x"FF",
x"FE",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"2C",
x"71",x"FF",x"FF",x"2C",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"71",x"FF",x"BA",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"FF",x"FA",x"F4",x"FF",x"FF",x"FF",x"FF",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F5",x"FF",x"FA",x"F4",
x"F4",x"F9",x"FF",x"FA",x"F4",x"F4",x"F4",x"FA",
x"FF",x"F5",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",
x"F5",x"FA",x"FF",x"F9",x"F4",x"F5",x"FA",x"FF",
x"FF",x"FF",x"F9",x"F4",x"F4",x"F5",x"FF",x"FF",
x"F4",x"F4",x"F4",x"F9",x"FF",x"FA",x"F4",x"FA",
x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"FA",x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",
x"FF",x"FF",x"FF",x"F5",x"F4",x"F4",x"F5",x"FF",
x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"96",x"FF",x"71",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"2C",x"FF",x"FF",x"2C",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F5",x"FF",
x"FF",x"F4",x"F4",x"FF",x"FF",x"FF",x"FA",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F9",x"FF",x"FA",x"F4",
x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",x"FA",x"FF",
x"F9",x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F5",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",
x"F5",x"F4",x"F4",x"F4",x"F4",x"FA",x"FF",x"F9",
x"F4",x"F4",x"F9",x"FF",x"FA",x"F4",x"F4",x"FE",
x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"FA",x"FF",x"F9",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",
x"FF",x"FF",x"FF",x"F4",x"F4",x"F4",x"F5",x"FF",
x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"B6",x"FF",x"4D",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"BA",x"FF",x"DB",
x"2C",x"8C",x"F4",x"F4",x"F4",x"FA",x"FF",x"FF",
x"F4",x"F4",x"F4",x"FF",x"FF",x"FF",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F9",x"FF",x"FA",x"F4",
x"F4",x"FF",x"FF",x"F5",x"F5",x"FF",x"FF",x"F9",
x"F4",x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",
x"F5",x"FA",x"FF",x"F9",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"FE",x"FF",x"F9",
x"F5",x"FE",x"FF",x"FE",x"F4",x"F4",x"F4",x"FE",
x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"FA",x"FF",x"FA",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",
x"FF",x"FF",x"FA",x"F4",x"F4",x"F4",x"F5",x"FF",
x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"2C",
x"96",x"FF",x"BA",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"2C",x"DB",x"FF",
x"FF",x"DA",x"FA",x"FE",x"FF",x"FF",x"FA",x"F4",
x"F4",x"F4",x"F4",x"FE",x"FF",x"FF",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F9",x"FF",x"FA",x"F4",
x"F4",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"F4",
x"F4",x"F4",x"F4",x"FF",x"FF",x"F5",x"F4",x"F4",
x"F4",x"FA",x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"FA",x"FF",x"FF",
x"FF",x"FF",x"FA",x"F4",x"F4",x"F4",x"F4",x"FA",
x"FF",x"FA",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F5",x"FF",x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FA",x"FF",x"F5",x"F4",x"F4",x"F4",
x"F9",x"FA",x"F4",x"F4",x"F4",x"F4",x"F9",x"FF",
x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F5",x"FF",x"FE",x"F9",x"DA",x"FF",
x"FF",x"BA",x"2C",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"71",
x"BA",x"FF",x"FF",x"FF",x"FA",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"FE",x"FF",x"F9",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F9",x"FF",x"FA",x"F4",
x"F4",x"F4",x"F9",x"FA",x"F5",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F5",x"F9",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F9",x"FA",
x"F9",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F9",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"FA",x"F9",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F9",x"FF",x"F5",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F9",x"FF",
x"FE",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FA",x"FF",x"FF",x"FF",x"FF",x"BA",
x"51",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F9",x"FA",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F9",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F5",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"90",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FF",x"F5",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FF",x"F9",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F9",x"FF",x"F9",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FA",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F5",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F9",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FF",x"F9",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FA",x"FA",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FF",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F5",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F5",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FF",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F5",x"F5",
x"F4",x"F4",x"F5",x"F9",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F5",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F5",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FF",x"FF",x"FF",x"FE",
x"F4",x"F4",x"F5",x"FF",x"F4",x"FA",x"FF",x"FF",
x"F4",x"F4",x"F4",x"FA",x"FE",x"FA",x"FF",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FA",x"FF",x"FF",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FF",x"F4",x"F4",x"F9",
x"F9",x"F4",x"F4",x"F4",x"F4",x"F4",x"FA",x"FA",
x"F4",x"F4",x"FF",x"FF",x"F4",x"F5",x"FF",x"F9",
x"F4",x"F4",x"FA",x"FE",x"F4",x"F4",x"F4",x"FA",
x"FF",x"FE",x"F9",x"F4",x"F4",x"F4",x"F9",x"FF",
x"FE",x"FA",x"F4",x"F4",x"F9",x"FF",x"F4",x"F4",
x"F4",x"F5",x"FA",x"F4",x"F4",x"F4",x"F4",x"FF",
x"F5",x"F4",x"F4",x"FA",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"FE",x"FA",x"F4",x"F9",x"FF",
x"F4",x"F4",x"F5",x"FF",x"F9",x"FA",x"F4",x"F9",
x"F4",x"F4",x"FA",x"FA",x"F4",x"FA",x"FA",x"F4",
x"F4",x"F4",x"F4",x"FA",x"FA",x"F4",x"FE",x"F5",
x"F4",x"F4",x"F5",x"FA",x"FF",x"FF",x"FF",x"FA",
x"F5",x"F4",x"F4",x"F4",x"F4",x"F4",x"FA",x"FE",
x"F4",x"FA",x"FA",x"FE",x"F5",x"FF",x"F9",x"FF",
x"F4",x"F4",x"F9",x"FF",x"F4",x"F4",x"FF",x"F9",
x"F4",x"F4",x"F4",x"F4",x"F4",x"FA",x"FA",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F5",x"FF",x"F4",x"F4",
x"F4",x"FF",x"FA",x"FF",x"F4",x"F4",x"F4",x"FF",
x"F5",x"F4",x"FF",x"FF",x"FA",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F9",x"FF",x"F4",x"F4",x"FF",x"FF",
x"F9",x"F4",x"F5",x"FF",x"FF",x"F4",x"F4",x"F4",
x"F4",x"F5",x"FF",x"FA",x"FF",x"F9",x"F4",x"F4",
x"F4",x"F4",x"FA",x"FE",x"F4",x"F4",x"FF",x"FA",
x"F5",x"FE",x"FA",x"F9",x"FF",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F9",x"FF",
x"F4",x"FF",x"F4",x"FE",x"FA",x"FF",x"F4",x"FF",
x"F4",x"F4",x"F9",x"FF",x"F4",x"F5",x"FF",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"FF",x"F5",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F5",x"FF",x"F4",x"F4",
x"FA",x"FF",x"F4",x"FA",x"FF",x"F4",x"F4",x"FF",
x"F9",x"F5",x"FA",x"F9",x"FE",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FF",x"F5",x"F4",x"F5",x"FA",x"FA",
x"FA",x"F4",x"F5",x"FF",x"FA",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FE",x"F5",x"F4",x"F4",x"F4",x"F9",
x"F4",x"F5",x"FF",x"F4",x"F4",x"FA",x"FF",x"FA",
x"F4",x"F4",x"F4",x"F4",x"FF",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F5",x"FF",
x"F9",x"FA",x"F4",x"FE",x"FF",x"F9",x"F4",x"FF",
x"F5",x"F4",x"F9",x"FF",x"F4",x"F4",x"FA",x"FF",
x"FE",x"FA",x"F4",x"F4",x"F4",x"F9",x"FF",x"FF",
x"FA",x"F5",x"F4",x"F4",x"F5",x"FF",x"F4",x"F4",
x"FF",x"F5",x"F4",x"F4",x"FA",x"FE",x"F4",x"FE",
x"F9",x"FE",x"F5",x"F5",x"FF",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F5",x"FF",x"F4",x"F4",x"FF",x"F4",x"F9",
x"FF",x"F4",x"F5",x"FF",x"F4",x"F4",x"F4",x"F4",
x"F4",x"FF",x"FA",x"F4",x"F4",x"F4",x"F9",x"FA",
x"F4",x"FF",x"F5",x"F4",x"F5",x"FF",x"FA",x"FA",
x"F4",x"F4",x"F4",x"F4",x"FF",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F5",x"FF",
x"FF",x"F5",x"F4",x"FE",x"FF",x"F4",x"F4",x"FE",
x"F9",x"F4",x"F5",x"FF",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F9",x"FF",x"FA",x"F4",x"F4",x"F4",x"F4",
x"F5",x"FA",x"FF",x"F4",x"F4",x"FF",x"F4",x"F4",
x"FF",x"F4",x"F4",x"F4",x"F9",x"FF",x"F4",x"FA",
x"FE",x"FF",x"F4",x"F9",x"FF",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F9",x"FE",x"F4",x"FF",x"F5",x"F4",x"F5",
x"FF",x"F4",x"F5",x"FF",x"F4",x"F4",x"F4",x"F4",
x"F4",x"FF",x"FA",x"F4",x"F4",x"F4",x"FF",x"F4",
x"F5",x"FF",x"F4",x"F4",x"FF",x"F5",x"FA",x"FA",
x"F4",x"F4",x"F4",x"F4",x"FF",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F5",x"FF",
x"FF",x"F4",x"F4",x"FF",x"FE",x"F4",x"F4",x"FE",
x"F9",x"F4",x"F5",x"FF",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"FF",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"FF",x"F4",x"F4",x"FF",x"F4",x"F5",
x"FF",x"F4",x"F4",x"F4",x"FF",x"FA",x"F4",x"FA",
x"FF",x"F9",x"F4",x"F9",x"FF",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F9",x"FF",x"FF",x"F9",x"F4",x"F4",x"F4",
x"FF",x"F4",x"F4",x"FF",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F9",x"FF",x"F9",x"F9",x"FF",x"F5",x"F4",
x"FA",x"FF",x"F9",x"FF",x"F5",x"F4",x"FA",x"FF",
x"F4",x"F4",x"F4",x"F4",x"FF",x"F5",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"FF",
x"FA",x"F4",x"F4",x"FF",x"F9",x"F4",x"F4",x"FE",
x"F9",x"F4",x"F4",x"FF",x"F4",x"F4",x"F4",x"F5",
x"F4",x"F4",x"FF",x"F9",x"F4",x"F4",x"F5",x"F4",
x"F4",x"FA",x"FE",x"F4",x"F4",x"FF",x"F4",x"F4",
x"FF",x"FA",x"F5",x"FF",x"FE",x"F4",x"F4",x"F9",
x"FF",x"F4",x"F4",x"FA",x"FF",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F5",x"F4",x"F4",x"F4",x"F4",x"F4",
x"FF",x"F4",x"F4",x"FF",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F5",x"FA",x"FA",x"F4",x"F4",x"F4",
x"F4",x"FA",x"FA",x"F4",x"F4",x"F4",x"F5",x"F9",
x"F4",x"F4",x"F4",x"F4",x"FA",x"F5",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"FF",
x"F4",x"F4",x"F4",x"F5",x"F4",x"F4",x"F4",x"FA",
x"F5",x"F4",x"F4",x"FF",x"F4",x"F4",x"F9",x"FF",
x"FF",x"FF",x"F9",x"F4",x"F4",x"F4",x"FF",x"FF",
x"FF",x"FA",x"F4",x"F4",x"F4",x"FF",x"F4",x"F4",
x"F5",x"FA",x"FA",x"F9",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"FA",x"FF",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F5",
x"FF",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"FA",
x"FE",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F9",x"FF",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F5",x"FE",x"FF",x"F5",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"FA",x"FA",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"8C",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"8C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E9",x"E9",x"E9",x"E4",x"E0",
x"E4",x"E9",x"E9",x"E9",x"E0",x"E0",x"E9",x"E9",
x"E9",x"E9",x"E0",x"E4",x"ED",x"E9",x"E0",x"E0",
x"E4",x"ED",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E9",x"E9",x"E0",x"E0",x"E4",x"E9",x"E9",x"E9",
x"E4",x"E4",x"E4",x"E0",x"E0",x"E9",x"E4",x"E9",
x"E9",x"E9",x"E9",x"E4",x"E9",x"E9",x"E9",x"E9",
x"E0",x"E9",x"E9",x"E9",x"E4",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"FF",x"F6",x"F6",x"FF",x"ED",
x"F6",x"F6",x"F2",x"F6",x"F6",x"E4",x"FF",x"F2",
x"F2",x"F2",x"E4",x"FB",x"F2",x"F6",x"F2",x"E9",
x"FB",x"F2",x"F6",x"ED",x"E0",x"E0",x"E4",x"FF",
x"F6",x"F2",x"FB",x"E4",x"F6",x"F6",x"F2",x"F2",
x"E9",x"F2",x"FF",x"E4",x"E0",x"FB",x"E9",x"F2",
x"F6",x"FB",x"F2",x"E9",x"FF",x"F2",x"F2",x"F2",
x"E0",x"FF",x"F2",x"F2",x"FB",x"ED",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"FF",x"ED",x"ED",x"FB",x"ED",
x"F6",x"F6",x"F2",x"F6",x"F6",x"E4",x"FF",x"F2",
x"F2",x"E0",x"E9",x"FF",x"F2",x"F2",x"E4",x"ED",
x"FB",x"F2",x"ED",x"E4",x"E0",x"E0",x"F2",x"F2",
x"E0",x"E0",x"E0",x"E0",x"F6",x"F6",x"F2",x"E9",
x"E0",x"F2",x"F6",x"FF",x"E4",x"FB",x"E4",x"E0",
x"ED",x"F2",x"E0",x"E0",x"FF",x"F2",x"F2",x"E0",
x"E0",x"FF",x"F2",x"F2",x"FB",x"ED",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"FF",x"F2",x"F2",x"ED",x"E0",
x"F6",x"F2",x"F2",x"FB",x"E0",x"E4",x"FF",x"E9",
x"E9",x"E0",x"E0",x"E9",x"ED",x"F2",x"FF",x"E0",
x"E9",x"ED",x"F6",x"FB",x"E0",x"E0",x"F2",x"F6",
x"E0",x"E0",x"E4",x"E0",x"F6",x"F2",x"E9",x"E4",
x"E0",x"F2",x"ED",x"E9",x"FF",x"FF",x"E4",x"E0",
x"ED",x"F2",x"E0",x"E0",x"FF",x"E9",x"E9",x"E0",
x"E0",x"FF",x"ED",x"F6",x"F6",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"FF",x"E4",x"E0",x"E0",x"E0",
x"F6",x"ED",x"E0",x"FB",x"F2",x"E4",x"FF",x"F6",
x"F6",x"F6",x"E9",x"FB",x"F6",x"FB",x"F6",x"E9",
x"FB",x"F6",x"FB",x"F2",x"E0",x"E0",x"E4",x"FB",
x"FB",x"F6",x"FB",x"E4",x"F6",x"FB",x"F6",x"F6",
x"ED",x"F2",x"ED",x"E0",x"E9",x"FF",x"E4",x"E0",
x"ED",x"F6",x"E0",x"E0",x"FF",x"F6",x"F6",x"F6",
x"E4",x"FF",x"E4",x"E0",x"FF",x"E9",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E4",x"E0",x"E0",x"E0",x"E0",
x"E4",x"E0",x"E0",x"E4",x"E4",x"E0",x"E4",x"E4",
x"E4",x"E4",x"E0",x"E0",x"E9",x"E4",x"E0",x"E0",
x"E0",x"E9",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E4",x"E4",x"E0",x"E0",x"E4",x"E4",x"E4",x"E4",
x"E4",x"E4",x"E0",x"E0",x"E0",x"E4",x"E0",x"E0",
x"E0",x"E4",x"E0",x"E0",x"E4",x"E4",x"E4",x"E4",
x"E0",x"E4",x"E0",x"E0",x"E4",x"E4",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"F6",
x"FB",x"FB",x"F6",x"E4",x"F2",x"ED",x"E0",x"E4",
x"F6",x"F2",x"FB",x"FB",x"FB",x"F6",x"FB",x"FB",
x"FB",x"FB",x"E9",x"E9",x"FB",x"FB",x"F2",x"E0",
x"E9",x"FB",x"E4",x"E0",x"ED",x"ED",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",
x"E9",x"E4",x"FB",x"ED",x"F6",x"ED",x"E0",x"E4",
x"FB",x"E0",x"E0",x"FF",x"E4",x"E0",x"E0",x"ED",
x"F2",x"E0",x"E9",x"FF",x"E4",x"E0",x"F6",x"F2",
x"E9",x"FF",x"FB",x"E0",x"F2",x"ED",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",
x"F6",x"F6",x"FB",x"E9",x"F6",x"ED",x"E0",x"E4",
x"FB",x"E0",x"E0",x"FF",x"E4",x"E0",x"E0",x"ED",
x"F2",x"E0",x"ED",x"F6",x"E0",x"E0",x"E9",x"FB",
x"E9",x"F6",x"F2",x"FB",x"F2",x"ED",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"FF",
x"E9",x"E4",x"F6",x"F2",x"F2",x"F6",x"E4",x"ED",
x"F6",x"E0",x"E0",x"FF",x"E4",x"E0",x"E0",x"ED",
x"F2",x"E0",x"E4",x"FF",x"E9",x"E4",x"FB",x"F2",
x"E9",x"F6",x"E0",x"F2",x"FF",x"ED",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"F2",
x"F6",x"F6",x"F2",x"E0",x"E4",x"F2",x"FB",x"F6",
x"E4",x"E0",x"E0",x"F2",x"E4",x"E0",x"E0",x"E9",
x"ED",x"E0",x"E0",x"E9",x"F6",x"F6",x"ED",x"E0",
x"E4",x"ED",x"E0",x"E0",x"F2",x"E9",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E4",x"E9",x"E9",x"E9",x"E9",
x"E0",x"E4",x"E9",x"E9",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E9",x"E9",x"E0",x"E4",x"E9",x"E9",x"E9",
x"E9",x"E0",x"E0",x"E9",x"E4",x"E0",x"E0",x"E9",
x"E9",x"E9",x"E4",x"E0",x"E9",x"E9",x"E9",x"E9",
x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E9",x"F2",x"FF",x"F6",x"F2",
x"E9",x"FF",x"F2",x"F6",x"FB",x"E0",x"E0",x"E0",
x"FB",x"F2",x"F2",x"FB",x"E9",x"F2",x"FB",x"F6",
x"F2",x"E0",x"E0",x"FF",x"F2",x"E0",x"E0",x"FB",
x"F6",x"F2",x"FB",x"F2",x"ED",x"F2",x"FF",x"F2",
x"E9",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"FB",x"E9",x"E0",
x"F6",x"ED",x"E0",x"E0",x"FB",x"ED",x"E0",x"E0",
x"FB",x"F6",x"F2",x"ED",x"E0",x"E0",x"F6",x"ED",
x"E0",x"E0",x"ED",x"F2",x"FF",x"E4",x"E0",x"FB",
x"F6",x"F2",x"FB",x"F2",x"E0",x"E4",x"FB",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"FB",x"E9",x"E0",
x"F6",x"ED",x"E0",x"E0",x"FB",x"E9",x"E0",x"E0",
x"E4",x"ED",x"ED",x"FF",x"E9",x"E0",x"F6",x"ED",
x"E0",x"E0",x"FF",x"F6",x"FF",x"F2",x"E0",x"FB",
x"ED",x"F2",x"FB",x"E0",x"E0",x"E4",x"FB",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"FB",x"E9",x"E0",
x"E4",x"FF",x"F6",x"FB",x"F6",x"E0",x"E0",x"E0",
x"FB",x"F6",x"F6",x"FF",x"E4",x"E0",x"F6",x"ED",
x"E0",x"ED",x"F2",x"E0",x"E0",x"FF",x"E4",x"FB",
x"E9",x"E0",x"FB",x"ED",x"E0",x"E4",x"FF",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E4",x"E0",x"E0",
x"E0",x"E0",x"E9",x"E4",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E4",x"E9",x"E0",x"E0",x"E0",x"E4",x"E0",
x"E0",x"E4",x"E0",x"E0",x"E0",x"E4",x"E0",x"E4",
x"E0",x"E0",x"E4",x"E4",x"E0",x"E0",x"E4",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"4C",x"91",x"91",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"4C",x"B5",x"91",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"4C",x"F9",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"B5",x"91",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"91",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"B5",x"4C",x"28",x"91",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"B5",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"4C",x"28",x"28",x"F9",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"4C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"91",x"91",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"91",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"4C",x"91",x"28",x"28",x"28",
x"28",x"28",x"91",x"91",x"28",x"28",x"28",x"4C",
x"F9",x"91",x"28",x"91",x"91",x"28",x"4C",x"91",
x"91",x"4C",x"28",x"4C",x"F9",x"91",x"28",x"F9",
x"91",x"91",x"28",x"28",x"91",x"91",x"28",x"28",
x"28",x"4C",x"91",x"4C",x"B5",x"B5",x"4C",x"91",
x"91",x"91",x"4C",x"91",x"91",x"4C",x"91",x"4C",
x"4C",x"28",x"4C",x"91",x"91",x"B5",x"91",x"4C",
x"28",x"4C",x"91",x"4C",x"4C",x"91",x"91",x"91",
x"91",x"91",x"91",x"91",x"28",x"28",x"91",x"91",
x"28",x"4C",x"91",x"4C",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"91",x"91",x"28",x"4C",x"91",
x"4C",x"B5",x"4C",x"28",x"B5",x"28",x"28",x"28",
x"F9",x"28",x"B5",x"4C",x"28",x"B5",x"28",x"F9",
x"91",x"28",x"28",x"28",x"F9",x"28",x"28",x"F9",
x"28",x"91",x"4C",x"B5",x"91",x"B5",x"91",x"28",
x"28",x"F9",x"28",x"4C",x"91",x"91",x"28",x"91",
x"B5",x"4C",x"28",x"28",x"B5",x"28",x"B5",x"4C",
x"91",x"91",x"4C",x"4C",x"91",x"91",x"28",x"F9",
x"4C",x"B5",x"91",x"F9",x"28",x"F9",x"91",x"28",
x"F9",x"91",x"28",x"F9",x"28",x"B5",x"91",x"B5",
x"91",x"F9",x"28",x"4C",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"B5",x"28",x"28",x"91",
x"28",x"F9",x"28",x"28",x"F9",x"28",x"28",x"28",
x"F9",x"28",x"F9",x"28",x"28",x"F9",x"28",x"F9",
x"28",x"28",x"28",x"28",x"F9",x"28",x"28",x"F9",
x"28",x"91",x"91",x"F9",x"28",x"28",x"28",x"28",
x"28",x"4C",x"B5",x"91",x"91",x"91",x"28",x"91",
x"91",x"28",x"B5",x"91",x"B5",x"28",x"4C",x"91",
x"91",x"B5",x"91",x"28",x"91",x"91",x"28",x"F9",
x"91",x"91",x"28",x"28",x"28",x"F9",x"28",x"28",
x"F9",x"28",x"28",x"F9",x"28",x"F9",x"28",x"28",
x"28",x"4C",x"B5",x"91",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"4C",x"B5",x"91",x"B5",
x"28",x"4C",x"B5",x"91",x"4C",x"28",x"28",x"4C",
x"F9",x"4C",x"4C",x"B5",x"91",x"4C",x"4C",x"F9",
x"4C",x"28",x"28",x"28",x"F9",x"91",x"4C",x"F9",
x"4C",x"B5",x"B5",x"4C",x"B5",x"91",x"4C",x"28",
x"28",x"B5",x"91",x"91",x"91",x"B5",x"4C",x"B5",
x"B5",x"28",x"B5",x"91",x"B5",x"4C",x"28",x"B5",
x"28",x"91",x"4C",x"28",x"91",x"B5",x"91",x"4C",
x"28",x"B5",x"91",x"91",x"4C",x"F9",x"4C",x"4C",
x"F9",x"4C",x"4C",x"F9",x"4C",x"4C",x"B5",x"91",
x"4C",x"B5",x"91",x"91",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"91",x"4C",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"4C",x"91",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"91",
x"4C",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"4C",x"F9",x"91",x"B5",x"4C",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"91",x"4C",x"4C",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"F9",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"F9",x"28",x"91",
x"91",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"F9",x"28",x"91",x"91",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"F9",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"B5",x"28",x"28",x"F9",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"91",
x"91",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"F9",x"91",x"91",x"4C",
x"4C",x"F9",x"28",x"B5",x"28",x"B5",x"B5",x"91",
x"91",x"28",x"28",x"28",x"91",x"B5",x"91",x"B5",
x"B5",x"28",x"B5",x"28",x"B5",x"4C",x"91",x"B5",
x"91",x"B5",x"B5",x"28",x"B5",x"4C",x"28",x"4C",
x"F9",x"91",x"B5",x"F9",x"B5",x"4C",x"B5",x"91",
x"4C",x"4C",x"F9",x"91",x"B5",x"91",x"B5",x"91",
x"28",x"28",x"4C",x"F9",x"91",x"28",x"F9",x"91",
x"B5",x"28",x"4C",x"91",x"B5",x"4C",x"28",x"28",
x"4C",x"91",x"F9",x"28",x"B5",x"B5",x"91",x"91",
x"B5",x"B5",x"28",x"B5",x"91",x"F9",x"28",x"91",
x"91",x"4C",x"B5",x"B5",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"F9",x"4C",x"B5",x"28",
x"28",x"F9",x"28",x"91",x"28",x"91",x"91",x"28",
x"F9",x"28",x"28",x"28",x"91",x"91",x"91",x"28",
x"F9",x"4C",x"B5",x"28",x"91",x"28",x"91",x"91",
x"91",x"28",x"F9",x"28",x"91",x"28",x"28",x"28",
x"F9",x"28",x"91",x"91",x"28",x"F9",x"28",x"28",
x"F9",x"28",x"F9",x"28",x"91",x"91",x"28",x"91",
x"28",x"28",x"28",x"F9",x"28",x"28",x"F9",x"28",
x"91",x"91",x"F9",x"91",x"91",x"4C",x"28",x"28",
x"4C",x"91",x"B5",x"28",x"91",x"91",x"28",x"F9",
x"28",x"F9",x"28",x"91",x"28",x"F9",x"28",x"91",
x"91",x"4C",x"B5",x"91",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"F9",x"28",x"91",x"B5",
x"28",x"F9",x"28",x"B5",x"28",x"91",x"91",x"28",
x"F9",x"28",x"28",x"91",x"91",x"28",x"91",x"28",
x"91",x"91",x"4C",x"F9",x"28",x"91",x"91",x"28",
x"91",x"28",x"91",x"B5",x"28",x"28",x"28",x"28",
x"F9",x"28",x"91",x"91",x"28",x"B5",x"4C",x"28",
x"B5",x"28",x"F9",x"28",x"91",x"91",x"28",x"91",
x"28",x"28",x"28",x"F9",x"28",x"28",x"F9",x"28",
x"91",x"91",x"B5",x"4C",x"28",x"28",x"28",x"28",
x"F9",x"28",x"91",x"28",x"91",x"91",x"28",x"F9",
x"28",x"91",x"F9",x"28",x"28",x"F9",x"28",x"91",
x"91",x"4C",x"28",x"B5",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"4C",x"91",x"4C",x"28",x"91",
x"4C",x"4C",x"91",x"4C",x"4C",x"91",x"91",x"4C",
x"91",x"4C",x"28",x"28",x"91",x"91",x"91",x"28",
x"28",x"4C",x"28",x"4C",x"28",x"28",x"91",x"91",
x"91",x"28",x"28",x"91",x"28",x"28",x"28",x"4C",
x"91",x"4C",x"91",x"91",x"28",x"28",x"91",x"91",
x"28",x"4C",x"91",x"4C",x"91",x"91",x"4C",x"91",
x"4C",x"28",x"28",x"91",x"91",x"4C",x"91",x"4C",
x"91",x"91",x"28",x"91",x"91",x"4C",x"28",x"28",
x"4C",x"91",x"91",x"4C",x"91",x"91",x"4C",x"91",
x"4C",x"28",x"4C",x"28",x"4C",x"91",x"4C",x"91",
x"91",x"4C",x"91",x"91",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"91",x"4C",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"4C",x"91",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0");
 
  constant ImageGO : GO_Screen := (
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",x"2C",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"C0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E4",x"ED",x"F2",
x"FB",x"FB",x"FF",x"FB",x"FB",x"F2",x"ED",x"E4",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E4",x"F2",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"F6",x"ED",x"E9",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E4",x"FB",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"F2",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E4",x"FB",x"FF",x"FF",x"FF",x"FF",x"F6",
x"ED",x"E4",x"E4",x"E4",x"E9",x"F2",x"FB",x"FF",
x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E9",x"E9",x"E9",x"E9",
x"E9",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E4",x"E9",x"E9",x"E9",x"E9",x"E9",x"E4",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E9",
x"E9",x"E9",x"E9",x"E9",x"E9",x"E0",x"E0",x"E4",
x"E9",x"E9",x"E9",x"E9",x"E9",x"E9",x"E9",x"E9",
x"E9",x"E9",x"E9",x"E9",x"E9",x"F2",x"E4",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"FB",x"FF",x"FF",x"FF",x"FF",x"E9",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"ED",
x"FF",x"F2",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"F2",x"FF",x"FF",x"FF",
x"FF",x"E9",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FF",x"FF",x"ED",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"F2",
x"FF",x"FF",x"FF",x"FF",x"ED",x"E0",x"E0",x"E4",
x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E9",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"ED",x"FF",x"FF",x"FF",x"FF",x"E9",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"ED",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",
x"FF",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F2",x"FF",x"FF",x"FF",x"FF",x"E9",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"F6",
x"FF",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"E9",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"F6",x"FF",x"FF",x"FF",x"F2",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"FB",x"FF",x"FF",x"FF",
x"FF",x"F2",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F2",x"FF",x"FF",x"FF",x"FF",x"FB",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E9",x"FF",
x"FF",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"F2",x"FF",x"FF",x"FF",x"ED",x"ED",x"ED",x"ED",
x"ED",x"ED",x"ED",x"ED",x"ED",x"F6",x"E9",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E4",
x"FF",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E9",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F2",x"FF",x"FF",x"FF",x"FF",x"FF",
x"ED",x"E0",x"E0",x"E0",x"E0",x"E0",x"F6",x"FF",
x"FF",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"F2",x"FF",x"FF",x"FB",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E4",
x"FF",x"FF",x"FF",x"FB",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FB",x"FF",x"FF",x"F2",x"FF",
x"FF",x"FF",x"F2",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F2",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FB",x"E0",x"E0",x"E0",x"E0",x"E9",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"F2",x"FF",x"FF",x"FB",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E9",
x"FF",x"FF",x"FF",x"FB",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F6",x"F6",x"F2",x"F2",x"F2",x"F2",
x"F2",x"F2",x"F2",x"F2",x"E4",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E9",x"FF",x"FF",x"FB",x"E0",x"F2",
x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F2",x"FF",x"FF",x"F6",x"FF",x"FF",
x"FF",x"ED",x"E0",x"E0",x"E0",x"FB",x"FF",x"FF",
x"F6",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"F2",x"FF",x"FF",x"FF",x"ED",x"ED",x"ED",x"ED",
x"ED",x"F2",x"F6",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E4",
x"FF",x"FF",x"FF",x"FB",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"F2",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FB",x"FF",x"FF",x"ED",x"E0",x"E4",
x"FF",x"FF",x"FF",x"F6",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F2",x"FF",x"FF",x"F6",x"ED",x"FF",
x"FF",x"FF",x"E4",x"E0",x"ED",x"FF",x"FF",x"F2",
x"ED",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"F2",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FB",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E4",
x"FB",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FB",x"FB",x"FB",x"FB",
x"FF",x"FF",x"FF",x"ED",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E9",x"FF",x"FF",x"FB",x"E0",x"E0",x"E0",
x"F2",x"FF",x"FF",x"FF",x"E9",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F2",x"FF",x"FF",x"F6",x"E0",x"FB",
x"FF",x"FF",x"F2",x"E4",x"FF",x"FF",x"FF",x"E4",
x"ED",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"F2",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FB",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"F6",x"FF",x"FF",x"FF",x"F2",x"E0",x"E0",x"E0",
x"E0",x"E0",x"ED",x"E4",x"E4",x"E4",x"E4",x"E4",
x"FB",x"FF",x"FF",x"ED",x"E0",x"E0",x"E0",x"E0",
x"E0",x"F6",x"FF",x"FF",x"FB",x"ED",x"ED",x"ED",
x"F2",x"FF",x"FF",x"FF",x"F6",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F2",x"FF",x"FF",x"F6",x"E0",x"E9",
x"FF",x"FF",x"FF",x"F6",x"FF",x"FF",x"ED",x"E0",
x"ED",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"F2",x"FF",x"FF",x"FB",x"E9",x"E4",x"E4",x"E4",
x"E4",x"E9",x"F2",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"ED",x"FF",x"FF",x"FF",x"FF",x"E9",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"FB",x"FF",x"FF",x"ED",x"E0",x"E0",x"E0",x"E0",
x"E9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"E9",x"E0",x"E0",
x"E0",x"E0",x"F2",x"FF",x"FF",x"F6",x"E0",x"E0",
x"F6",x"FF",x"FF",x"FF",x"FF",x"FB",x"E0",x"E0",
x"ED",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"F2",x"FF",x"FF",x"FB",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"F6",x"FF",x"FF",x"FF",x"FF",x"ED",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E9",
x"FF",x"FF",x"FF",x"ED",x"E0",x"E0",x"E0",x"E0",
x"F6",x"FF",x"FF",x"F6",x"F2",x"F2",x"F2",x"F2",
x"F2",x"F6",x"FF",x"FF",x"FF",x"FB",x"E0",x"E0",
x"E0",x"E0",x"F2",x"FF",x"FF",x"F6",x"E0",x"E0",
x"E9",x"FF",x"FF",x"FF",x"FF",x"E9",x"E0",x"E0",
x"ED",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"F2",x"FF",x"FF",x"FB",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E4",x"FB",x"FF",x"FF",x"FF",x"FF",x"FB",
x"F2",x"E9",x"E9",x"E9",x"ED",x"F2",x"FB",x"FF",
x"FF",x"FF",x"FF",x"FB",x"E4",x"E0",x"E0",x"E9",
x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"E9",x"E0",
x"E0",x"E0",x"F2",x"FF",x"FF",x"F6",x"E0",x"E0",
x"E0",x"F6",x"FF",x"FF",x"F6",x"E0",x"E0",x"E0",
x"ED",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"F2",x"FF",x"FF",x"FB",x"E9",x"E9",x"E9",x"E9",
x"E9",x"E9",x"E9",x"E9",x"E9",x"ED",x"F2",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E4",x"FB",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"F6",x"E9",x"E0",x"E0",x"E0",x"F6",
x"FF",x"FF",x"F2",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"FB",x"E0",
x"E0",x"E0",x"F2",x"FF",x"FF",x"F6",x"E0",x"E0",
x"E0",x"E4",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"ED",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F2",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"ED",x"FB",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",
x"F6",x"E9",x"E0",x"E0",x"E0",x"E0",x"ED",x"FF",
x"FF",x"FF",x"F2",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E4",x"FB",x"FF",x"FF",x"FF",x"F2",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FB",x"E4",x"E0",
x"E0",x"E0",x"F2",x"F2",x"E0",x"E0",x"E0",x"E0",
x"F2",x"FF",x"FF",x"FF",x"ED",x"E0",x"E0",x"E0",
x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F2",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E4",x"E9",x"F2",
x"F6",x"FB",x"FB",x"F6",x"F6",x"ED",x"E9",x"E4",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"ED",x"ED",
x"ED",x"ED",x"E9",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E4",x"ED",x"ED",x"ED",x"ED",x"ED",
x"E4",x"E4",x"ED",x"ED",x"ED",x"ED",x"E4",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E9",x"ED",x"ED",x"ED",x"E9",x"E0",x"E0",x"E4",
x"ED",x"ED",x"ED",x"ED",x"ED",x"ED",x"ED",x"ED",
x"ED",x"ED",x"ED",x"ED",x"ED",x"F2",x"F2",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E4",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E4",x"E9",x"ED",x"ED",x"ED",x"E9",
x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E4",
x"E4",x"E4",x"E4",x"E4",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E4",x"E4",x"E4",x"E4",x"E4",
x"E0",x"E0",x"E4",x"E4",x"E4",x"E4",x"E4",x"E4",
x"E4",x"E4",x"E4",x"E4",x"E4",x"E4",x"E4",x"ED",
x"E4",x"E0",x"E0",x"E4",x"E4",x"E4",x"E4",x"E4",
x"E4",x"E4",x"E4",x"E4",x"E4",x"E4",x"E4",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E9",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FB",x"F2",x"E4",x"E0",x"E0",x"E0",x"E0",x"F6",
x"FF",x"FF",x"FF",x"FB",x"E9",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E4",x"FB",x"FF",x"FF",x"FF",x"F6",
x"E0",x"E4",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"E4",x"E0",x"E0",x"F6",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FB",
x"ED",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E4",x"F6",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"E9",x"E0",x"E0",x"E0",x"E4",
x"FF",x"FF",x"FF",x"FF",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"F2",x"FF",x"FF",x"FF",x"E4",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"E4",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"F6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"F6",x"FF",
x"FF",x"FF",x"FF",x"F2",x"ED",x"E9",x"ED",x"FB",
x"FF",x"FF",x"FF",x"FF",x"E9",x"E0",x"E0",x"E0",
x"F2",x"FF",x"FF",x"FF",x"E9",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"FF",x"FF",x"FF",x"F2",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FF",x"F2",x"F2",
x"F2",x"F2",x"F2",x"F2",x"F2",x"F2",x"F2",x"FB",
x"E4",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"F6",
x"F2",x"F2",x"F2",x"F2",x"F2",x"F6",x"FF",x"FF",
x"FF",x"FF",x"E9",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"ED",x"FF",x"FF",
x"FF",x"FB",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",
x"ED",x"FF",x"FF",x"FF",x"FB",x"E4",x"E0",x"E0",
x"E4",x"FF",x"FF",x"FF",x"F6",x"E0",x"E0",x"E0",
x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"E4",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FB",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E4",
x"E0",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"E4",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E9",x"FF",
x"FF",x"FF",x"F2",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"FB",x"FF",x"FF",
x"FB",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"F2",x"FF",x"FF",x"FF",x"ED",x"E0",x"E0",
x"E0",x"F2",x"FF",x"FF",x"FF",x"E9",x"E0",x"E0",
x"E0",x"E0",x"FB",x"FF",x"FF",x"F6",x"E0",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FB",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"E4",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E4",x"FF",
x"FF",x"FF",x"F2",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E9",x"FF",x"FF",x"FF",
x"F2",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E4",x"FF",x"FF",x"FF",x"F6",x"E0",x"E0",
x"E0",x"E4",x"FF",x"FF",x"FF",x"F6",x"E0",x"E0",
x"E0",x"ED",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FF",x"E9",x"E9",
x"E9",x"E9",x"E9",x"E9",x"F2",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"E9",
x"E4",x"E4",x"E4",x"E4",x"E4",x"E9",x"F6",x"FF",
x"FF",x"FF",x"ED",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E9",x"FF",x"FF",x"FF",
x"E9",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FB",x"FF",x"FF",x"FB",x"E0",x"E0",
x"E0",x"E0",x"F2",x"FF",x"FF",x"FF",x"E4",x"E0",
x"E0",x"FB",x"FF",x"FF",x"F6",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"F6",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FB",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",
x"E9",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FB",x"E0",x"E0",
x"E0",x"E0",x"E4",x"FF",x"FF",x"FF",x"F2",x"E0",
x"E9",x"FF",x"FF",x"FF",x"E4",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"F6",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"F6",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E9",x"FF",x"FF",x"FF",
x"ED",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"FB",x"FF",x"FF",x"FB",x"E0",x"E0",
x"E0",x"E0",x"E0",x"F6",x"FF",x"FF",x"FF",x"E4",
x"F6",x"FF",x"FF",x"F6",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FF",x"ED",x"ED",
x"ED",x"ED",x"ED",x"ED",x"F2",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"F2",
x"F2",x"F2",x"F6",x"FF",x"FF",x"FF",x"FB",x"E4",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E4",x"FF",x"FF",x"FF",
x"F6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E9",x"FF",x"FF",x"FF",x"F2",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E4",x"FF",x"FF",x"FF",x"F6",
x"FF",x"FF",x"FF",x"E9",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FB",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E4",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"E4",
x"E0",x"E0",x"E0",x"F6",x"FF",x"FF",x"FF",x"E9",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"F6",x"FF",x"FF",
x"FF",x"ED",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E4",x"FB",x"FF",x"FF",x"FF",x"E9",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"F6",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FB",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FB",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"E4",
x"E0",x"E0",x"E0",x"E4",x"FB",x"FF",x"FF",x"FB",
x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E4",x"FF",x"FF",
x"FF",x"FF",x"F2",x"E4",x"E0",x"E0",x"E0",x"E9",
x"FB",x"FF",x"FF",x"FF",x"F6",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E9",x"FF",x"FF",x"FF",
x"FF",x"FF",x"E9",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FB",x"E4",x"E4",
x"E4",x"E4",x"E4",x"E4",x"E4",x"E4",x"E4",x"E4",
x"ED",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"E4",
x"E0",x"E0",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",
x"F6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"ED",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FB",x"FB",x"FF",x"FF",
x"FF",x"FF",x"FF",x"F6",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"F6",x"FF",x"FF",
x"FF",x"FB",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"F2",x"E0",x"E0",x"ED",x"FF",x"FF",x"FF",x"E4",
x"E0",x"E0",x"E0",x"E0",x"E0",x"F2",x"FF",x"FF",
x"FF",x"ED",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E9",
x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"F2",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"F2",x"FF",x"FF",
x"FF",x"F6",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F6",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"F2",x"E0",x"E0",x"F2",x"FF",x"FF",x"FF",x"E9",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E9",x"FF",x"FF",
x"FF",x"FF",x"E9",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E9",x"F2",x"FB",x"FF",x"FF",x"FB",x"F6",
x"ED",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E4",x"F2",x"F2",x"F2",
x"F2",x"F2",x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E4",x"F2",x"F2",x"F2",x"F2",x"F2",x"F2",
x"F2",x"F2",x"F2",x"F2",x"F2",x"F2",x"F2",x"F6",
x"F2",x"E0",x"E4",x"F2",x"F2",x"F2",x"F2",x"ED",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E9",x"F2",x"F2",
x"F2",x"F2",x"F2",x"E4",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E4",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"64",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"2C",x"4C",x"4C",x"2C",x"28",x"2C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"6C",x"B0",x"6C",x"B0",x"4C",x"B0",x"2C",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"6C",x"90",x"28",x"6C",x"6C",x"B0",x"2C",
x"4C",x"90",x"90",x"4C",x"4C",x"90",x"90",x"6C",
x"4C",x"90",x"90",x"6C",x"2C",x"90",x"90",x"90",
x"2C",x"28",x"2C",x"90",x"90",x"90",x"2C",x"6C",
x"90",x"90",x"4C",x"4C",x"90",x"90",x"6C",x"28",
x"28",x"6C",x"4C",x"2C",x"8C",x"4C",x"B0",x"B0",
x"4C",x"4C",x"6C",x"28",x"90",x"2C",x"90",x"B0",
x"6C",x"28",x"2C",x"90",x"90",x"90",x"28",x"8C",
x"90",x"90",x"2C",x"8C",x"90",x"90",x"2C",x"90",
x"B0",x"6C",x"6C",x"90",x"90",x"2C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"6C",x"B0",x"8C",x"B0",x"4C",x"B0",x"4C",
x"B0",x"6C",x"6C",x"90",x"4C",x"4C",x"6C",x"B0",
x"6C",x"B0",x"4C",x"4C",x"4C",x"B0",x"4C",x"B0",
x"4C",x"28",x"2C",x"B0",x"4C",x"4C",x"4C",x"B0",
x"6C",x"6C",x"90",x"90",x"90",x"6C",x"B0",x"2C",
x"28",x"4C",x"B0",x"6C",x"6C",x"B0",x"4C",x"2C",
x"B0",x"4C",x"90",x"28",x"B0",x"2C",x"B0",x"6C",
x"28",x"28",x"2C",x"D0",x"4C",x"4C",x"4C",x"B0",
x"2C",x"6C",x"4C",x"B0",x"2C",x"90",x"6C",x"B0",
x"6C",x"4C",x"B0",x"6C",x"90",x"6C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"6C",x"90",x"2C",x"2C",x"28",x"B0",x"4C",
x"B0",x"6C",x"4C",x"4C",x"90",x"90",x"6C",x"B0",
x"2C",x"6C",x"90",x"B0",x"6C",x"B0",x"4C",x"4C",
x"2C",x"28",x"28",x"4C",x"8C",x"B0",x"6C",x"B0",
x"6C",x"4C",x"4C",x"B0",x"6C",x"4C",x"4C",x"2C",
x"28",x"2C",x"B0",x"B0",x"4C",x"B0",x"4C",x"2C",
x"D0",x"4C",x"90",x"28",x"B0",x"2C",x"B0",x"4C",
x"28",x"28",x"28",x"4C",x"90",x"B0",x"6C",x"B0",
x"28",x"4C",x"6C",x"90",x"28",x"6C",x"6C",x"B0",
x"4C",x"4C",x"B0",x"4C",x"4C",x"4C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"6C",x"90",x"28",x"28",x"28",x"B0",x"2C",
x"90",x"6C",x"90",x"6C",x"90",x"6C",x"90",x"B0",
x"6C",x"90",x"6C",x"B0",x"4C",x"B0",x"6C",x"B0",
x"4C",x"28",x"2C",x"B0",x"6C",x"B0",x"6C",x"90",
x"6C",x"90",x"6C",x"6C",x"90",x"6C",x"90",x"28",
x"28",x"28",x"6C",x"B0",x"28",x"6C",x"90",x"8C",
x"90",x"2C",x"B0",x"6C",x"D0",x"2C",x"B0",x"4C",
x"28",x"28",x"4C",x"B0",x"4C",x"B0",x"4C",x"B0",
x"6C",x"B0",x"4C",x"B0",x"6C",x"B0",x"4C",x"B0",
x"4C",x"2C",x"B0",x"6C",x"90",x"4C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"2C",x"2C",x"28",x"28",x"28",x"2C",x"28",
x"2C",x"4C",x"4C",x"2C",x"2C",x"4C",x"4C",x"2C",
x"2C",x"4C",x"4C",x"2C",x"28",x"2C",x"4C",x"2C",
x"28",x"28",x"28",x"2C",x"4C",x"4C",x"28",x"2C",
x"4C",x"4C",x"28",x"28",x"4C",x"4C",x"2C",x"28",
x"28",x"2C",x"6C",x"6C",x"28",x"2C",x"4C",x"4C",
x"2C",x"28",x"4C",x"4C",x"4C",x"28",x"2C",x"2C",
x"28",x"28",x"28",x"4C",x"4C",x"4C",x"28",x"2C",
x"4C",x"2C",x"28",x"2C",x"4C",x"4C",x"28",x"2C",
x"2C",x"28",x"2C",x"4C",x"4C",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"4C",x"6C",x"2C",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"4C",x"4C",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"6C",x"2C",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"6C",x"2C",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"4C",x"28",x"4C",x"4C",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"4C",x"8C",
x"28",x"2C",x"6C",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"4C",x"90",x"90",x"4C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"6C",x"90",x"4C",x"2C",x"28",x"2C",x"4C",
x"4C",x"28",x"B0",x"4C",x"2C",x"4C",x"4C",x"2C",
x"4C",x"2C",x"2C",x"2C",x"2C",x"2C",x"28",x"28",
x"4C",x"2C",x"2C",x"4C",x"4C",x"2C",x"28",x"28",
x"4C",x"B0",x"4C",x"6C",x"90",x"4C",x"2C",x"28",
x"2C",x"4C",x"4C",x"28",x"28",x"28",x"6C",x"D0",
x"6C",x"2C",x"B0",x"28",x"2C",x"4C",x"4C",x"28",
x"4C",x"28",x"4C",x"4C",x"2C",x"28",x"4C",x"2C",
x"4C",x"4C",x"28",x"8C",x"4C",x"4C",x"B0",x"2C",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"6C",x"B0",x"6C",x"B0",x"2C",x"B0",x"6C",
x"B0",x"4C",x"B0",x"4C",x"90",x"6C",x"90",x"6C",
x"90",x"4C",x"B0",x"6C",x"90",x"4C",x"28",x"28",
x"90",x"4C",x"90",x"90",x"8C",x"6C",x"28",x"28",
x"4C",x"B0",x"4C",x"6C",x"B0",x"6C",x"B0",x"2C",
x"90",x"6C",x"90",x"6C",x"28",x"28",x"6C",x"90",
x"B0",x"2C",x"B0",x"2C",x"B0",x"6C",x"B0",x"4C",
x"B0",x"6C",x"90",x"8C",x"6C",x"4C",x"8C",x"B0",
x"6C",x"90",x"2C",x"28",x"4C",x"8C",x"90",x"2C",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"6C",x"8C",x"28",x"B0",x"6C",x"B0",x"8C",
x"90",x"6C",x"B0",x"4C",x"B0",x"2C",x"4C",x"B0",
x"6C",x"B0",x"B0",x"90",x"90",x"2C",x"28",x"28",
x"B0",x"4C",x"B0",x"4C",x"4C",x"90",x"28",x"28",
x"2C",x"B0",x"2C",x"6C",x"90",x"2C",x"B0",x"4C",
x"D0",x"6C",x"90",x"8C",x"28",x"28",x"6C",x"6C",
x"6C",x"90",x"B0",x"4C",x"D0",x"6C",x"90",x"6C",
x"4C",x"D0",x"4C",x"4C",x"B0",x"90",x"4C",x"B0",
x"90",x"6C",x"2C",x"28",x"4C",x"6C",x"B0",x"2C",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"6C",x"90",x"2C",x"B0",x"6C",x"B0",x"2C",
x"4C",x"4C",x"B0",x"4C",x"B0",x"4C",x"4C",x"90",
x"4C",x"D0",x"8C",x"B0",x"90",x"28",x"28",x"28",
x"B0",x"4C",x"90",x"4C",x"4C",x"90",x"28",x"28",
x"2C",x"B0",x"2C",x"6C",x"8C",x"2C",x"B0",x"4C",
x"B0",x"2C",x"4C",x"4C",x"28",x"28",x"6C",x"6C",
x"2C",x"B0",x"B0",x"4C",x"B0",x"2C",x"4C",x"4C",
x"6C",x"B0",x"8C",x"28",x"B0",x"B0",x"2C",x"6C",
x"2C",x"B0",x"6C",x"6C",x"2C",x"2C",x"D0",x"2C",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"4C",x"90",x"90",x"8C",x"2C",x"8C",x"90",
x"90",x"2C",x"90",x"2C",x"6C",x"90",x"90",x"4C",
x"28",x"90",x"4C",x"6C",x"4C",x"28",x"28",x"28",
x"8C",x"4C",x"6C",x"4C",x"4C",x"6C",x"28",x"28",
x"2C",x"90",x"6C",x"4C",x"6C",x"2C",x"90",x"2C",
x"6C",x"90",x"90",x"4C",x"28",x"28",x"4C",x"6C",
x"28",x"4C",x"90",x"28",x"8C",x"90",x"90",x"2C",
x"90",x"2C",x"90",x"2C",x"8C",x"6C",x"28",x"90",
x"90",x"90",x"4C",x"6C",x"90",x"90",x"6C",x"2C",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"2C",x"2C",x"28",x"28",x"28",x"2C",
x"2C",x"28",x"2C",x"28",x"28",x"2C",x"2C",x"28",
x"28",x"2C",x"28",x"28",x"28",x"28",x"28",x"28",
x"2C",x"28",x"2C",x"28",x"28",x"2C",x"28",x"28",
x"28",x"2C",x"2C",x"28",x"28",x"28",x"2C",x"28",
x"28",x"2C",x"2C",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"2C",x"28",x"28",x"2C",x"2C",x"28",
x"2C",x"28",x"2C",x"4C",x"B0",x"2C",x"28",x"28",
x"2C",x"2C",x"28",x"28",x"2C",x"2C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"2C",x"2C",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"2C",x"2C",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"2C",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"6C",x"6C",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"4C",x"90",x"2C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"6C",x"B0",x"90",x"6C",x"28",x"6C",x"90",
x"6C",x"2C",x"6C",x"90",x"90",x"4C",x"4C",x"90",
x"6C",x"4C",x"90",x"90",x"B0",x"2C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"6C",x"90",x"2C",x"B0",x"4C",x"B0",x"2C",
x"90",x"6C",x"6C",x"4C",x"90",x"6C",x"4C",x"B0",
x"4C",x"90",x"6C",x"4C",x"B0",x"2C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"6C",x"8C",x"28",x"B0",x"6C",x"90",x"28",
x"6C",x"90",x"90",x"8C",x"90",x"90",x"4C",x"90",
x"28",x"B0",x"4C",x"4C",x"B0",x"2C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"6C",x"B0",x"4C",x"B0",x"4C",x"B0",x"4C",
x"B0",x"6C",x"B0",x"4C",x"90",x"90",x"4C",x"90",
x"28",x"90",x"6C",x"6C",x"B0",x"2C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"2C",x"4C",x"6C",x"4C",x"28",x"4C",x"6C",
x"4C",x"2C",x"4C",x"6C",x"4C",x"4C",x"2C",x"4C",
x"28",x"2C",x"6C",x"6C",x"4C",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"2C",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"2C",x"28",x"28",x"28",
x"28",x"2C",x"4D",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"71",
x"4C",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"71",x"BA",x"B6",x"2C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"2C",x"71",x"2C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"2C",x"2C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"2C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"2C",
x"2C",x"2C",x"2C",x"4D",x"DB",x"96",x"96",x"B6",
x"96",x"71",x"DB",x"2C",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"2C",x"DB",
x"71",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"2C",x"DF",x"4D",x"96",x"96",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"4D",x"DF",x"4D",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"2C",x"96",x"71",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"51",x"96",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"51",
x"BA",x"BA",x"BA",x"B6",x"FF",x"96",x"51",x"51",
x"51",x"51",x"DB",x"2C",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"2C",x"DB",
x"71",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"95",x"BA",x"28",x"2C",x"4D",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"4D",x"DB",x"2C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"2C",x"2C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"96",x"BA",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"2C",
x"4D",x"2C",x"28",x"28",x"FF",x"4D",x"28",x"28",
x"28",x"4D",x"DB",x"2C",x"28",x"71",x"B6",x"4D",
x"28",x"28",x"28",x"28",x"2C",x"71",x"51",x"28",
x"2C",x"4D",x"28",x"28",x"2C",x"2C",x"2C",x"DB",
x"71",x"28",x"28",x"2C",x"2C",x"2C",x"2C",x"4D",
x"96",x"71",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"BA",x"95",x"28",x"28",x"28",x"28",x"2C",
x"2C",x"28",x"28",x"2C",x"4D",x"2C",x"51",x"96",
x"2C",x"28",x"28",x"28",x"28",x"4C",x"51",x"2C",
x"28",x"28",x"28",x"28",x"4D",x"DB",x"2C",x"28",
x"28",x"28",x"2C",x"71",x"4D",x"28",x"2C",x"2C",
x"28",x"28",x"4D",x"2C",x"4D",x"71",x"28",x"4D",
x"4D",x"28",x"2C",x"2C",x"28",x"28",x"28",x"2C",
x"71",x"96",x"4D",x"2C",x"28",x"96",x"96",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"FF",x"51",x"28",x"28",
x"28",x"4C",x"DB",x"2C",x"4D",x"DA",x"96",x"B6",
x"28",x"28",x"28",x"4D",x"BA",x"96",x"DB",x"2C",
x"51",x"DB",x"2C",x"51",x"DB",x"71",x"28",x"BA",
x"71",x"2C",x"51",x"BA",x"DB",x"71",x"96",x"BA",
x"71",x"51",x"28",x"28",x"28",x"28",x"28",x"28",
x"2C",x"BA",x"96",x"51",x"71",x"4D",x"51",x"DB",
x"71",x"2C",x"28",x"4D",x"DF",x"71",x"BA",x"BA",
x"71",x"28",x"28",x"28",x"28",x"96",x"FF",x"BA",
x"96",x"4D",x"2C",x"28",x"4D",x"DB",x"2C",x"28",
x"28",x"51",x"BA",x"96",x"BA",x"2C",x"B6",x"51",
x"28",x"28",x"DA",x"71",x"71",x"DA",x"28",x"96",
x"96",x"2C",x"96",x"DB",x"2C",x"28",x"2C",x"96",
x"BA",x"96",x"FF",x"4D",x"28",x"96",x"96",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"DF",x"51",x"28",x"28",
x"28",x"2C",x"DB",x"2C",x"BA",x"71",x"51",x"BA",
x"2C",x"28",x"2C",x"BA",x"71",x"2C",x"DB",x"4D",
x"4D",x"DB",x"4D",x"BA",x"96",x"96",x"28",x"BA",
x"96",x"96",x"BA",x"4D",x"2C",x"71",x"DB",x"2C",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"71",
x"BA",x"FF",x"BA",x"96",x"95",x"4D",x"DB",x"96",
x"DB",x"BA",x"2C",x"4D",x"FF",x"DB",x"4C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"DB",x"51",
x"51",x"96",x"96",x"2C",x"4D",x"DB",x"2C",x"28",
x"4D",x"DB",x"51",x"4D",x"DB",x"2C",x"B6",x"71",
x"28",x"2C",x"DB",x"51",x"71",x"DB",x"28",x"96",
x"BA",x"4D",x"BA",x"BA",x"71",x"28",x"71",x"BA",
x"2C",x"71",x"FF",x"71",x"28",x"96",x"96",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"DF",x"51",x"28",x"28",
x"28",x"2C",x"DB",x"71",x"BA",x"2C",x"4D",x"DB",
x"2C",x"2C",x"B6",x"96",x"2C",x"96",x"FF",x"51",
x"4C",x"DB",x"95",x"96",x"71",x"BA",x"28",x"BA",
x"FF",x"96",x"2C",x"28",x"28",x"4D",x"BA",x"B6",
x"71",x"4D",x"2C",x"28",x"28",x"28",x"28",x"2C",
x"2C",x"BA",x"71",x"28",x"28",x"4D",x"FF",x"2C",
x"2C",x"BA",x"96",x"4D",x"FF",x"96",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"DB",x"4D",
x"28",x"28",x"96",x"96",x"51",x"DB",x"2C",x"2C",
x"BA",x"71",x"2C",x"B6",x"FF",x"4D",x"71",x"B6",
x"28",x"51",x"FF",x"4D",x"51",x"DB",x"28",x"71",
x"BA",x"96",x"71",x"BA",x"71",x"2C",x"DB",x"51",
x"2C",x"BA",x"BA",x"96",x"28",x"96",x"96",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"DF",x"51",x"28",x"28",
x"28",x"2C",x"DB",x"DB",x"71",x"28",x"4D",x"DB",
x"2C",x"71",x"DB",x"2C",x"51",x"BA",x"DB",x"51",
x"2C",x"DB",x"DB",x"4D",x"71",x"BA",x"2C",x"BA",
x"DB",x"2C",x"28",x"28",x"28",x"28",x"28",x"4D",
x"71",x"BA",x"B6",x"28",x"28",x"28",x"28",x"28",
x"28",x"B6",x"96",x"28",x"28",x"71",x"BA",x"28",
x"28",x"71",x"BA",x"4D",x"FF",x"2C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"2C",x"DB",x"51",
x"2C",x"4D",x"BA",x"71",x"51",x"DB",x"2C",x"71",
x"BA",x"2C",x"71",x"BA",x"DB",x"4D",x"4D",x"DB",
x"4D",x"BA",x"FF",x"4C",x"51",x"DB",x"28",x"51",
x"FF",x"BA",x"2C",x"BA",x"71",x"51",x"DB",x"2C",
x"96",x"71",x"71",x"BA",x"28",x"71",x"96",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"FF",x"51",x"28",x"28",
x"28",x"2C",x"FF",x"DF",x"2C",x"28",x"4D",x"DB",
x"2C",x"BA",x"75",x"4D",x"BA",x"4D",x"DB",x"71",
x"2C",x"DB",x"DA",x"2C",x"71",x"BA",x"28",x"96",
x"FF",x"BA",x"96",x"4D",x"2C",x"28",x"28",x"2C",
x"28",x"4D",x"DB",x"28",x"28",x"28",x"28",x"28",
x"28",x"96",x"96",x"28",x"28",x"96",x"BA",x"2C",
x"2C",x"DB",x"71",x"2C",x"FF",x"2C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"96",x"FF",x"BA",
x"B6",x"96",x"71",x"2C",x"51",x"DB",x"2C",x"DB",
x"71",x"51",x"BA",x"4D",x"DB",x"4D",x"2C",x"96",
x"DB",x"BA",x"DB",x"2C",x"4D",x"DB",x"2C",x"4D",
x"FF",x"95",x"2C",x"BA",x"71",x"96",x"BA",x"96",
x"B6",x"2C",x"4D",x"FF",x"28",x"2C",x"2C",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"DF",x"4D",x"28",x"28",
x"28",x"28",x"FF",x"96",x"28",x"28",x"51",x"DB",
x"2C",x"BA",x"DB",x"DA",x"51",x"28",x"BA",x"71",
x"28",x"96",x"71",x"28",x"96",x"BA",x"28",x"71",
x"DB",x"2C",x"96",x"DB",x"B6",x"4D",x"71",x"96",
x"96",x"DA",x"51",x"28",x"28",x"28",x"28",x"28",
x"28",x"96",x"96",x"28",x"28",x"4D",x"DF",x"B6",
x"DB",x"96",x"28",x"2C",x"FF",x"2C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"2C",x"DB",x"51",
x"28",x"28",x"28",x"28",x"4D",x"DB",x"4D",x"DB",
x"BA",x"BA",x"4D",x"2C",x"DB",x"51",x"28",x"2C",
x"2C",x"51",x"DB",x"2C",x"4D",x"DB",x"2C",x"2C",
x"96",x"2C",x"2C",x"DB",x"71",x"51",x"DB",x"96",
x"2C",x"28",x"2C",x"FF",x"2C",x"51",x"BA",x"2C",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"2C",x"28",x"28",x"28",
x"28",x"28",x"B6",x"4D",x"28",x"28",x"4C",x"96",
x"2C",x"2C",x"4D",x"2C",x"28",x"28",x"2C",x"2C",
x"28",x"28",x"28",x"28",x"51",x"71",x"28",x"2C",
x"71",x"28",x"28",x"28",x"28",x"2C",x"71",x"96",
x"71",x"2C",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"96",x"96",x"28",x"28",x"28",x"2C",x"4D",
x"2C",x"28",x"28",x"28",x"51",x"2C",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"DB",x"4D",
x"28",x"28",x"28",x"28",x"28",x"2C",x"28",x"2C",
x"4D",x"2C",x"28",x"28",x"2C",x"2C",x"28",x"28",
x"28",x"71",x"DB",x"28",x"2C",x"51",x"2C",x"28",
x"28",x"28",x"2C",x"71",x"4D",x"28",x"28",x"28",
x"28",x"28",x"4C",x"FF",x"2C",x"2C",x"71",x"2C",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"51",x"71",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"DB",x"51",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"71",x"DB",x"2C",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"96",x"BA",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"96",x"4D",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"28",x"4D",x"BA",x"2C",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"2C",x"71",x"DF",x"51",x"28",x"28",x"28",x"28",
x"28",x"28",x"28",x"28",x"28",x"28",x"28",x"28",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"BA",x"FF",x"D5",x"90",x"90",x"90",x"90",x"90",
x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"90",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F9",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",
x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4",x"F4");
  constant kokoro : kokoroImage := ( 
 x"00",x"00",x"6D",x"6D",x"6D",x"6D",x"00",x"00",
x"00",x"00",x"6D",x"6D",x"6D",x"6D",x"00",x"00",
x"00",x"6D",x"C0",x"C0",x"C0",x"6D",x"6D",x"00",
x"00",x"6D",x"6D",x"C0",x"C0",x"C0",x"6D",x"00",
x"6D",x"C0",x"C0",x"C0",x"C0",x"C0",x"6D",x"6D",
x"6D",x"6D",x"C0",x"C0",x"C0",x"C0",x"C0",x"6D",
x"6D",x"C0",x"C0",x"FF",x"FF",x"C0",x"C0",x"6D",
x"6D",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"6D",
x"6D",x"C0",x"C0",x"FF",x"FF",x"C0",x"C0",x"C0",
x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"6D",
x"6D",x"C0",x"FF",x"FF",x"FF",x"C0",x"C0",x"C0",
x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"6D",
x"6D",x"C0",x"FF",x"FF",x"C0",x"C0",x"C0",x"C0",
x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"6D",
x"6D",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",
x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"6D",
x"00",x"6D",x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",
x"C0",x"C0",x"C0",x"C0",x"C0",x"C0",x"6D",x"00",
x"00",x"00",x"6D",x"C0",x"C0",x"C0",x"C0",x"C0",
x"C0",x"C0",x"C0",x"C0",x"C0",x"6D",x"00",x"00",
x"00",x"00",x"00",x"6D",x"C0",x"C0",x"C0",x"C0",
x"C0",x"C0",x"C0",x"C0",x"6D",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"6D",x"C0",x"C0",x"C0",
x"C0",x"C0",x"C0",x"6D",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"6D",x"C0",x"C0",x"C0",
x"C0",x"C0",x"C0",x"6D",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"6D",x"C0",x"C0",
x"C0",x"C0",x"6D",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"6D",x"C0",
x"C0",x"6D",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6D",
x"6D",x"00",x"00",x"00",x"00",x"00",x"00",x"00");
  
  constant duck : characterImage := (
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"00",x"00",x"00",x"00",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"00",
x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"FF",
x"00",x"00",x"00",x"00",x"FF",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"FF",x"FF",x"FF",x"FF",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"00",x"00",x"00",
x"00",x"00",x"00",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"D0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"D0",x"D0",
x"D0",x"D0",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"4D",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"4D",x"4D",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"4D",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"FF",
x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4D",
x"4D",x"4D",x"4D",x"4D",x"4D",x"4D",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"92",x"FF",x"FF",x"FF",
x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4D",
x"4D",x"4D",x"4D",x"4D",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"92",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"4D",x"4D",x"4D",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"92",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"4D",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"92",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"92",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"D0",x"D0",x"D0",x"D0",x"D0",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"92",x"92",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"D0",x"D0",x"D0",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"92",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"D0",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"92",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"92",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"92",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"92",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"92",x"92",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"92",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"92",x"92",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"92",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"92",x"92",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"92",x"92",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"92",x"92",x"92",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"92",x"92",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"92",x"92",
x"92",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"92",x"92",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"92",x"92",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"92",x"92",x"92",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"92",x"92",x"92",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"92",
x"92",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"92",x"92",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"92",x"92",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"92",
x"92",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"D0",x"D0",x"D0",x"D0",x"D0",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"D0",x"D0",x"D0",x"D0",x"D0",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"D0",x"D0",x"D0",x"D0",x"D0",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"D0",x"D0",x"D0",x"D0",x"D0",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"D0",x"D0",x"D0",x"D0",x"D0",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"D0",x"D0",x"D0",x"D0",x"D0",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"D0",x"D0",x"D0",
x"D0",x"00",x"00",x"D0",x"D0",x"D0",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"D0",x"D0",x"D0",x"D0",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"D0",x"D0",
x"D0",x"D0",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"D0",x"D0",x"D0",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"D0",x"D0",x"00",x"00",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"D0",x"D0",x"00",x"00",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"D0",x"D0",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"D0",x"D0",x"D0",x"00",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"D0",x"D0",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"D0",
x"D0",x"D0",x"D0",x"00",x"00",x"00",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"D0",x"D0",x"D0",x"D0",
x"D0",x"00",x"00",x"00",x"00",x"00",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"D0",x"D0",x"D0",x"D0",x"D0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"D0",x"D0",x"D0",x"D0",x"D0",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"D0",x"D0",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"D0",x"D0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");
constant strawberry : objectImage := (
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"55",x"55",x"55",x"55",x"E0",x"E0",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"55",x"55",x"55",x"E0",x"E0",x"E0",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"55",x"55",x"E0",x"E0",x"E0",x"E0",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"E0",x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"E0",x"E0",
x"E0",x"E0",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"F8",x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"F8",
x"F8",x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"E0",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"F8",
x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"55",x"55",x"55",x"55",x"55",x"55",
x"55",x"55",x"E0",x"E0",x"E0",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"55",x"55",x"55",x"55",x"55",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"55",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"55",
x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"E0",
x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"F8",x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"E0",
x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"F8",x"F8",x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"E0",
x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"F8",x"F8",x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"55",x"E0",x"E0",
x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"F8",x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"55",x"E0",x"E0",x"E0",
x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"55",x"E0",x"E0",x"E0",x"E0",
x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",x"55",
x"55",x"55",x"55",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"F8",x"F8",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",x"55",
x"55",x"55",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",x"F8",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",
x"55",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",x"F8",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F8",x"F8",x"F8",x"F8",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"55",x"55",x"55",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F8",x"F8",x"F8",x"F8",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F8",x"F8",x"F8",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"F8",
x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",x"E0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"F8",x"F8",
x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",x"E0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",x"F8",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",
x"F8",x"E0",x"E0",x"E0",x"E0",x"E0",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",
x"E0",x"E0",x"E0",x"E0",x"E0",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"F8",x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"F8",x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"F8",x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"F8",x"F8",x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"F8",x"F8",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",x"E0",
x"E0",x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",
x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",x"F8",x"E0",
x"E0",x"E0",x"E0",x"E0",x"F8",x"F8",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"E0",x"E0",
x"E0",x"E0",x"E0",x"F8",x"F8",x"F8",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",
x"E0",x"E0",x"E0",x"F8",x"F8",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",x"E0",
x"E0",x"E0",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"E0",x"E0",x"E0",x"E0",
x"E0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");
constant Anviel : objectImage := (
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"49",
x"49",x"49",x"49",x"49",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"49",
x"49",x"49",x"49",x"49",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"49",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"49",
x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"00",
x"00",x"00",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"49",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"49",
x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",
x"92",x"92",x"92",x"92",x"92",x"92",x"00",x"00",
x"00",x"00",x"00",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"49",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"49",
x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",
x"92",x"92",x"92",x"92",x"92",x"00",x"00",x"00",
x"00",x"00",x"00",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"49",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"49",
x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",
x"49",x"92",x"92",x"92",x"92",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"49",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"49",
x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",
x"49",x"92",x"92",x"92",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"49",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"49",
x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",
x"49",x"49",x"49",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"92",
x"92",x"92",x"92",x"92",x"49",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",
x"49",x"49",x"49",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",
x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"49",x"49",x"49",x"24",
x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",
x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",
x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"92",x"92",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",
x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",
x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"49",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");

	
  
 -- signal next_state, present_state : State_Values;  
	--Embbeded signals
	--For moving an object in the x axis
  signal xButton  : integer range 0 to 640;
   --For making objects fall 
  signal yButton  : integer range 0 to 500;
  signal yButton2 : integer range 0 to 500;
  
  --Offsets of all objects in screen
  signal offsetXP  : STD_LOGIC_VECTOR (9 downto 0);
  signal offsetYP  : STD_LOGIC_VECTOR (9 downto 0);
  signal offsetXF  : STD_LOGIC_VECTOR (9 downto 0);
  signal offsetYF  : STD_LOGIC_VECTOR (9 downto 0);
  signal offsetXA  : STD_LOGIC_VECTOR (9 downto 0);
  signal offsetYA  : STD_LOGIC_VECTOR (9 downto 0);
  signal offsetXC  : STD_LOGIC_VECTOR (9 downto 0);
  signal offsetYC  : STD_LOGIC_VECTOR (9 downto 0);
  signal offsetXGO : STD_LOGIC_VECTOR (9 downto 0) := "0010000000";--fixed offset
  signal offsetYGO : STD_LOGIC_VECTOR (9 downto 0) := "0010110000";--fixed offset
  
  signal offsetXBS : STD_LOGIC_VECTOR (9 downto 0) := "0010000000";--fixed offset
  signal offsetYBS : STD_LOGIC_VECTOR (9 downto 0) := "0010110000";--fixed offset
  
  --Addresses that are used for making large operations
  signal SuperAddressP : STD_LOGIC_VECTOR (16 downto 0);
  signal SuperAddressC : STD_LOGIC_VECTOR (13 downto 0);
  signal SuperAddressF : STD_LOGIC_VECTOR (15 downto 0);
  signal SuperAddressA : STD_LOGIC_VECTOR (15 downto 0);
  signal SuperAddressGO: STD_LOGIC_VECTOR (16 downto 0);
  signal SuperAddressBS: STD_LOGIC_VECTOR (16 downto 0);


  --For knowing when an element is touched by the duck
  signal flag          : STD_LOGIC;
  signal flagA         : STD_LOGIC;
  --Toggle for when the duck just touched the strawberry
  signal flagScore     : STD_LOGIC;
  --Toggle for when the duck just touched the anviel
  signal FlagHeart     : STD_LOGIC;
  signal FlagOutH      : STD_LOGIC;
  signal extraOffsetXC : STD_LOGIC_VECTOR(5 downto 0);
  --Signal that helps first draw and then remove hearts
  signal hearties : integer range 0 to 48;
  --Toggle for when the start button is pressed
  signal startFlag     : STD_LOGIC;
  
  
begin

   --Calculates the address that will be taken from the memory for each object
  SuperAddressP <= (Xin-offsetXP) + ((Yin-offsetYP)&"0000000");
  AddressChar <= SuperAddressP(13 downto 0);
  
  SuperAddressC <= (Xin-offsetXC - extraOffsetXC) + ((Yin-offsetYC)&"0000");
  AddressKok <= SuperAddressC(7 downto 0);

  SuperAddressF <= (Xin-offsetXF) + ((Yin - offsetYF)&"000000");
  AddressObj <= SuperAddressF(11 downto 0);
  
  SuperAddressA <= (Xin-offsetXA) + ((Yin - offsetYA)&"000000");
  AddressObj2 <= SuperAddressA(11 downto 0);
  
  SuperAddressGO <= (Xin-offsetXGO) + ((Yin - offsetYGO)&"0000000");
  AddressGO <= SuperAddressGO(13 downto 0);
  
  SuperAddressBS <= (Xin-offsetXBS) + ((Yin - offsetYBS)&"0000000");
  AddressBS <= SuperAddressBS(13 downto 0);
  
  Start_Screen: process (rst) 
  begin
		if(rst = '1')then
			startFlag <= '1';
		else 
			startFlag <= '0';
		end if; 
  end process Start_Screen;
  
  
  Corazon: process (enable2 , rst , clk)
  begin
    -- Check if pixel is in the active zone
	 if (rst = '1') then 
		 hearties <= 48;   --Pixels shown
		 offsetYC <= "0001010000";
		 offsetXC <= "0000110000";
	 elsif(rising_edge(clk)) then		
-- if the anviel crashes with the duck, one heart is removed by restricting the drawing zone for the hearts	 
		if(flagoutH = '1' and hearties /= 0) then
			hearties <= hearties - 16;  -- Reducing the number of pixels equivalent of one heart
		end if;
	 end if;
  end process Corazon;
  
  ExtraOffset: process(rst, clk)
  begin
		if (rst = '1')then
			extraOffsetXC <= "000000";
		elsif(rising_edge(Clk)) then
			if((Xin-offsetXC) >= 32) then
				extraOffsetXC <= "100000";
			elsif((Xin-offsetXC) >= 16) then 
				extraOffsetXC <= "010000";
			else
				extraOffsetXC <= "000000";
			end if;
		end if;
		
  end process ExtraOffset;
  
 --The next process updates the duck's positions according to the inputs from buttons
  Pato: process (rightB, leftB, enable60,rst, xButton, clk)
  begin
	 if (rst = '1') then
		--Initial values (places duck in the middle)
		 xbutton <= 256;
		 offsetYP <= "0101100000";
		 offsetXP <= CONV_STD_LOGIC_VECTOR(512, 10);
	 elsif(rising_edge(clk)) then
		if(enable60 = '1') then
		 -- Updates the offset in Y 
			offsetXP <= CONV_STD_LOGIC_VECTOR(640 - xButton, 10);
			if (rightB = '1' and xbutton > 0) then
			-- If clicked to the right, the value of the button decreases
				xButton <= xButton - 1;
			elsif (leftB = '1' and xbutton < 512) then
			-- If clicked to the left, the value of the button increases
				xButton <= xButton + 1;
			end if;
		end if;
	 end if;
  end process Pato;
  
  
 --The next process updates the strawberrie's positions according to the inputs from buttons
  Fresa: process (rightB, leftB, enable2 ,rst, yButton, clk)
  begin
	 if (rst = '1') then
			--Initial values 
		 ybutton <= 0;
		 offsetYF <= "0000000000";
		 offsetXF <= CONV_STD_LOGIC_VECTOR(288, 10); 
	 elsif(rising_edge(clk)) then
		if(Enable2 = '1') then
		   -- Makes the offset increase, so it goes down the screen
			yButton <= yButton + 1;
		elsif(yButton = 480) then
		   offsetXF <= offsetXF + 64; 
			yButton <= 0;
		end if;
		offsetYF <= CONV_STD_LOGIC_VECTOR(yButton, 10);
	 end if;
  end process Fresa;
   
	
	
	--The next process updates the anviel's positions according to the inputs from buttons
    Yunque: process (rightB, leftB, enable3, rst, yButton2, clk)
  begin
	 if (rst = '1') then
		-- Initial values
		 ybutton2 <= 0;
		 offsetYA <= "0000000000";
		 offsetXA <= CONV_STD_LOGIC_VECTOR(520, 10);
	 elsif(rising_edge(clk)) then
		if(yButton2 = 480) then
			offsetXA <= offsetXP - 64;
			yButton2 <= 0;
		elsif(Enable3= '1') then
		   -- Makes Y offset increase, so it goes down the screen
			yButton2 <= yButton2 + 1;
		end if;
		offsetYA <= CONV_STD_LOGIC_VECTOR(yButton2, 10);
	 end if;
  end process Yunque;

  
  process (En,Xin, Yin, addressChar, xButton, offsetYF, offsetYA, flag, addressObj, offsetXA, offsetXF, offsetXC, offsetYC) 
  begin
--	if(rst = '1')then
--		startFlag <= '1';
--	else 
--		startFlag <= '0';
--	end if; 
    -- Check if pixel is in the active zone
		if (En = '1') then
		--Checks if the reset or start button is pressed
			if (startFlag = '0') then
			
				if (Xin >= 256 and Xin < 384 and Yin >= 176 and Yin < 304) then
					Color <= ImageBS (conv_integer(AddressBS));
				else 
					Color <="00000000";
				end if;
				
			elsif(hearties = 0) then
				if (Xin >= 256 and Xin < 384 and Yin >= 176 and Yin < 304) then
					Color <= ImageGO (conv_integer(AddressGO));
				else 
					Color <="00000000";
				end if;
			
			elsif ((Xin >= offsetXC and Xin < (offsetXC + hearties) and Yin >= offsetYC and Yin < offsetYC + 16)
			and kokoro(conv_integer(AddressKok)) /= "00000000") then
			 
				Color <= kokoro (conv_integer(AddressKok));
			
			--For drawing the strawberry, we must check:
			 -- *If the Xin and Yin are in the place the strawberry will be drawn
			 -- *If the color that will be drawn is not black
			 -- *If it has not been touched by the duck
			 elsif ( (Xin>= offsetXF and Xin < (offsetXF + 64)) and Yin >= offsetYF and Yin < 64 + offsetYF and 
			 strawberry(conv_integer(AddressObj)) /= "00000000" and flag = '0') then
				  
					Color <= strawberry(conv_integer(AddressObj));
			
			--For drawing the anviel, we must check:
			 -- *If the Xin and Yin are in the place the anviel will be drawn
			 -- *If the color that will be drawn is not black
			 -- *If it has not been touched by the duck
			  elsif ( (Xin>= offsetXA and Xin < (offsetXA + 64)) and Yin >= offsetYA and Yin < 64 + offsetYA and 
			  Anviel(conv_integer(AddressObj2)) /= "00000000"  and flagA = '0') then
				  
						Color <= Anviel(conv_integer(AddressObj2));
			--For drawing the duck, we must check if the Xin and Yin are in the place the duck will be drawn
			  elsif ((Xin>= (512 - xButton) and Xin < (640 - xButton)) and Yin > 352) then
				 Color <= duck (conv_integer(AddressChar));
			  else
				 --In any other case, draw everything black
				 Color <= "00000000"; -- Black
			  end if;
	 else
			-- EXTREMLY IMPORTANT
			-- Not in active zone, pixels should be OFF
			Color <= "00000000"; -- Off
	 end if;
  end process;


	--The next process checks if the duck touches the strawberry
  CollisionCheck: process (offsetYF, offsetYP, offsetXP, offsetXF, flag) 
  begin
	if(rising_edge(clk)) then
		--First, check if the middle from the bottom line of the stawbeerry is inside the space of the duck
		if ((offsetYF + 46) > offsetYP and offsetXP > (offsetXF + 32) and (offsetXP - 128) < (offsetXF + 32)
		and (offsetYF + 64) < 480) then
			flag <= '1';
		--Second, check if the duck has alraedy touched the strawberry and the it is below the Y offset of the duck
		elsif (flag = '1' and (offsetYF + 64) > offsetYP and (offsetYF) < 480) then
			flag <= '1';
		else 
		--In any other case, it is 0. The strawberry must be drawn
			flag <= '0';
		end if;
	end if;
  end process CollisionCheck;
  
  
  
  --The next process checks if the duck touches the anviel
  CrashCheck: process (offsetYA, offsetYP, offsetXP, offsetXA, flagA)
  begin
	if(rising_edge(clk)) then
		--First, check if the middle from the bottom line of the anviel is inside the space of the duck
			if ((offsetYA + 46) > offsetYP and offsetXP > (offsetXA + 32) and (offsetXP - 128) < (offsetXA + 32) 
			and (offsetYA + 64) < 480) then
				flagA <= '1';
		--Second, check if the duck has alraedy touched the anviel and the it is below the Y offset of the duck
			elsif (flagA = '1' and (offsetYA + 64) > offsetYP and (offsetYA) < 480) then
				flagA <= '1';
			else 
		--In any other case, it is 0. The anviel must be drawn
				flagA <= '0';
			end if;
	 end if;
  end process CrashCheck;
  
  --The next process sends a one pulse 
  ScoreCheck: process(rst, clk, flagScore, flag)
  begin
   if (rst = '1') then
		flagScore <= '0';
		flagOut <= '0';
	elsif (rising_edge(Clk)) then 
		if (flagScore = '0' and flag = '1') then
			flagScore <= '1';
			FlagOut <= '1';
		elsif (flagscore = '1' and (offsetYF + 64) > offsetYP) then
			flagScore <= '1';
			FlagOut <= '0';
		else 
			flagScore <= '0';
			FlagOut <= '0';
		end if;
	end if;
  end process ScoreCheck;
  
 -- This process together with the CrashCheck one helps us remove hearts (lifes)
  HeartOff: process(rst, clk, flagHeart, flagA)
  begin
   if (rst = '1') then
		FlagHeart <= '0';
		FlagOutH <= '0';
	elsif (rising_edge(Clk)) then 
		if (flagHeart = '0' and flagA = '1') then
			flagHeart <= '1';
			flagOutH  <= '1';
		elsif (flagHeart = '1' and (offsetYA + 64) > offsetYP) then
			FlagHeart <= '1';
			flagOutH  <= '0';
		else 
			FlagOutH  <= '0';
			FlagHeart <= '0';
		end if;
	end if;
  end process HeartOff;

  -- Send individual color to their channel
  R <= Color(7 downto 5);
  G <= Color(4 downto 2);
  B <= Color(1 downto 0);

end Behavioral;





